// serial_out.v

// Generated using ACDS version 23.1 993
`default_nettype none
module serial_out (
    input wire clk,          // System clock
    input wire reset_n,      // Active-low reset
    input wire uart_tx       // UART TX line (connected to your module)
	);

    wire [7:0] rx_data;       // Data received from UART
    wire rx_valid;            // UART data valid flag
    reg [31:0] av_writedata;  // Data to write to JTAG UART
    reg av_write_n;           // Write signal for JTAG UART (active low)
    wire av_waitrequest;      // Waitrequest signal from JTAG UART

    // Avalon-MM signals for the JTAG UART
    reg av_chipselect;        // Chip select for JTAG UART
    reg av_address;     // Address for JTAG UART
    reg av_read_n;            // Read signal (not used in this example)
    wire [31:0] av_readdata;  // Read data (not used in this example)
    wire av_irq;              // Interrupt request (not used in this example)
	wire readyfordata;

    reg [7:0] temp_data = 8'd65;

    // Instantiate UART Receiver
    uart_rx uart_rx_inst (
        .clk(clk),
        .reset_n(reset_n),
        .rx(uart_tx),
        .data(rx_data),
        .valid(rx_valid)
    );

	// // Handle the writing of data to the JTAG UART
    // always @(posedge clk or negedge reset_n) begin
    //     if (!reset_n) begin
    //         av_writedata <= {24'b0, temp_data};
    //         av_write_n <= 1'b0; // Disabled by default
    //         av_chipselect <= 1'b1;
    //         av_address <= 1'b0;
    //         av_read_n <= 1'b1;
    //         temp_data <= 8'd65;
    //     end else begin
    //         av_writedata <= {24'b0, temp_data}; // Write 8-bit UART data to JTAG UART (32-bit word)
    //         av_write_n <= 1'b0;               // Active low, so write when 0
    //         av_chipselect <= 1'b1;            // Enable chip select to JTAG UART
    //         av_address <= 1'b0;            // Address for data register (depends on your design)
    //         av_read_n <= 1'b1;
	// 		   if (!av_waitrequest && readyfordata) begin
    //             if(temp_data >= 8'd90) begin
    //                 temp_data <= 8'd65;
    //             end
    //             else begin
    //                 temp_data <= temp_data + 1;
    //             end
	// 		   end
	// 			else begin
	// 			    temp_data <= temp_data;
	// 			end
    //     end
    // end

    // Handle the writing of data to the JTAG UART
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            av_writedata <= 0;
            av_write_n <= 1'b1; // Disabled by default
            av_chipselect <= 0;
            av_address <= 0;
            av_read_n <= 1'b1;
        end else if (rx_valid) begin
            av_writedata <= {24'b0, rx_data}; // Write 8-bit UART data to JTAG UART (32-bit word)
            av_write_n <= 1'b0;               // Active low, so write when 0
            av_chipselect <= 1'b1;            // Enable chip select to JTAG UART
            av_address <= 1'b0;            // Address for data register (depends on your design)
        end 
		  else if (!av_waitrequest && readyfordata) begin
            av_write_n <= 1'b1;               // No write if JTAG UART is not ready
            av_chipselect <= 0;               // Disable chip select
        end
    end

    // Instantiate JTAG UART
	serial_out_jtag_uart_0 jtag_uart_0_kavish (
		.clk            (clk), //               clk.clk
		.rst_n          (reset_n), //             reset.reset_n
		.av_chipselect  (av_chipselect), // avalon_jtag_slave.chipselect
		.av_address     (av_address), //                  .address
		.av_read_n      (av_read_n), //                  .read_n
		.av_readdata    (av_readdata), //                  .readdata
		.av_write_n     (av_write_n), //                  .write_n
		.av_writedata   (av_writedata), //                  .writedata
		.av_waitrequest  (av_waitrequest), //                  .waitrequest
		.av_irq         (av_irq),  //               irq.irq
		.readyfordata   (readyfordata)
	);

endmodule


