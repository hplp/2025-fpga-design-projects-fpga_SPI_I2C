
module serial_out (
	);	

endmodule
