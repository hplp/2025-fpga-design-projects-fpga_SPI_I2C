	component serial_out is
	end component serial_out;

	u0 : component serial_out
		port map (
		);

