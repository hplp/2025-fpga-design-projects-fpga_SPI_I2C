`default_nettype none
module servive
(
 input wire 	   i_clk,
 input wire 	   i_rst_n,
 output wire 	   q,
 output wire 	   uart_txd);

   parameter memfile = "zephyr_hello.hex";
   parameter memsize = 8192;

   wire      wb_clk;
   wire      wb_rst;

   assign uart_txd = q;

   servive_clock_gen clock_gen
     (.i_clk (i_clk),
      .i_rst (!i_rst_n),
      .o_clk (wb_clk),
      .o_rst (wb_rst));

   servant_spi_top
     #(.memfile (memfile),
       .memsize (memsize))
   servant
     (.wb_clk (wb_clk),
      .wb_rst (wb_rst),
      .q      (q));
		
	serial_out serial_out
		(.clk(i_clk),
       .reset_n(i_rst_n),
       .uart_tx(q));

endmodule
